typedef struct packed {
    logic [4:0] rs1;
    logic [4:0] rs2;
    logic [4:0] rd;
    logic en_rs1;
    logic en_rs2;
    logic en_rd;
    logic [63:0] immed;
    logic keep_pc_plus_immed;
    logic alu_use_immed;
    logic alu_width_32;
    logic [2:0] funct3;
    logic [6:0] funct7;
    logic is_store;
    logic is_load;
    logic is_csr;
    logic csr_rw;
    logic csr_rs;
    logic csr_rc;
    logic csr_immed;
    logic is_ecall;
    logic is_break;
    logic is_trap_ret;
    logic is_wfi;
    logic is_sfence_vma;
    logic is_atomic;
    logic alu_op;
    logic is_swap;
    logic alu_nop;
} decoder_output;
